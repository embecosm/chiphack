
module edge_detect(
  /* Here we need to input our buttons and the clock
      And to output the edge detect signal
  */
  );

  // The buttons on the mystorm are "active low" (they read as 1 when not pressed, and 0 when pressed)

  // We then have to produce a slower clock

  // Then we follow Saar's edge detect tutorial, but using the slow clock  

endmodule
