
module basics(

//////////// CLOCK //////////
input 		          		CLOCK_50,
//////////// LED //////////
output		     [7:0]		LED,
//////////// KEY //////////
input 		     [1:0]		KEY,
//////////// SW //////////
input 		     [3:0]		SW,
//////////// SDRAM //////////
output		    [12:0]		DRAM_ADDR,
output		     [1:0]		DRAM_BA,
output		          		DRAM_CAS_N,
output		          		DRAM_CKE,
output		          		DRAM_CLK,
output		          		DRAM_CS_N,
inout 		    [15:0]		DRAM_DQ,
output		     [1:0]		DRAM_DQM,
output		          		DRAM_RAS_N,
output		          		DRAM_WE_N,
//////////// EPCS //////////
output		          		EPCS_ASDO,
input 		          		EPCS_DATA0,
output		          		EPCS_DCLK,
output		          		EPCS_NCSO,
//////////// Accelerometer and EEPROM //////////
output		          		G_SENSOR_CS_N,
input 		          		G_SENSOR_INT,
output		          		I2C_SCLK,
inout 		          		I2C_SDAT,
//////////// ADC //////////
output		          		ADC_CS_N,
output		          		ADC_SADDR,
output		          		ADC_SCLK,
input 		          		ADC_SDAT,
//////////// 2x13 GPIO Header //////////
inout 		    [12:0]		GPIO_2,
input 		     [2:0]		GPIO_2_IN

);


/*
Register instantiation
*/
reg  [31:00] count;
reg          a;
reg          b;

/*
Wire instantiation
*/
wire [07:00] led_out;

/*
An 'assign' statement is simply connecting wires together, 
either directly or through logic
*/

// assign the most significant bit of the counter to be
// the LEd clock
assign led_clock = count[15];

// the edge detect signal is (b AND (NOT a))
assign ed = b & !a;

// connect the edge detect signal to an LED
assign led_out = {count[31:24]};
assign LED[07:00] = led_out;
// or
// assign LED[7:0] = count[15:08] 


// assign meaningful names to pushbutton keys
assign reset = KEY[0];
assign button = KEY[1];

/*
All synchronous logic need a clock, and most typically we
want the logic to change on the positive edge of the clock
*/

// simple counter to divide up the clock in order
// to create a slower frequency clock
always @(posedge CLOCK_50) begin
  if (reset == 1'b0) begin
    count <= 0;
  end
  else begin
    count <= count + 1;
    /* all the following statements are equivalent:
    count[15:00] <= count[15:0] + 1;
    count <= count + 1'b1;
    count <= count + 16'b0000000000000001;
    count[15:0] <= count + 16'h0001
    */
  end
end

always @(posedge led_clock) begin
  // it's always good to have a reset condition, otherwise
  // the state of the register will show up as undertemined
  // in simulation ('x')
  if (reset == 1'b0) begin
    a <= 0;
    b <= 0;	 
  end
  else begin
    // the pushbutton wire input is connected to the input
    // of a register / flip flop
    a <= button;
    b <= a;
  end
end


endmodule
