module mem #(parameter ABITS=9) (
	input clk,
	input [ABITS-1:0] addr,
	input [15:0] d,
	input rd,
	input wr,
	output reg [15:0] q,
	output wait
);

//`define testwithdelay 1
	reg [15:0] m[0:(1<<ABITS)-1];
	wire rdenable = rd & ~wait;
	wire wrenable = wr & ~wait;
	always @(posedge clk) begin
		if (rdenable)
			q <= m[addr];
		if (wrenable)
			m[addr] <= d;
	end

`ifndef testwithdelay
	assign wait = 0;
`else
	reg [1:0] delay;
	assign wait = delay != 2'd3;
	always @(posedge clk)
	if (~(rd|wr))
		delay <= 0;
	else if (delay != 2'd3)
		delay <= delay + 1;
`endif

	initial begin
/* initial orders */
		m[0]  <= (("T"-"@")<<11) | 30;
		m[1]  <= (("T"-"@")<<11) | 32;
		m[2]  <= (("T"-"@")<<11) | 31;
		m[3]  <= (("I"-"@")<<11) | 0;
		m[4]  <= (("S"-"@")<<11) | 33;
		m[5]  <= (("G"-"@")<<11) | 3;
		m[6]  <= (("L"-"@")<<11) | 11;
		m[7]  <= (("T"-"@")<<11) | 30;
		m[8]  <= (("I"-"@")<<11) | 0;
		m[9]  <= (("S"-"@")<<11) | 34;
		m[10] <= (("G"-"@")<<11) | 8;
		m[11] <= (("T"-"@")<<11) | 32;
		m[12] <= (("A"-"@")<<11) | 31;
		m[13] <= (("V"-"@")<<11) | 35;
		m[14] <= (("L"-"@")<<11) | 16;
		m[15] <= (("A"-"@")<<11) | 32;
		m[16] <= (("T"-"@")<<11) | 31;
		m[17] <= (("I"-"@")<<11) | 0;
		m[18] <= (("S"-"@")<<11) | 34;
		m[19] <= (("E"-"@")<<11) | 11;
		m[20] <= (("T"-"@")<<11) | 0;
		m[21] <= (("A"-"@")<<11) | 31;
		m[22] <= (("A"-"@")<<11) | 30;
		m[23] <= (("T"-"@")<<11) | 37;
		m[24] <= (("A"-"@")<<11) | 23;
		m[25] <= (("A"-"@")<<11) | 36;
		m[26] <= (("U"-"@")<<11) | 23;
		m[27] <= (("S"-"@")<<11) | 37;
		m[28] <= (("G"-"@")<<11) | 1;
		m[29] <= (("E"-"@")<<11) | 37;
		m[30] <= (("@"-"@")<<11) | 0;
		m[31] <= (("@"-"@")<<11) | 0;
		m[32] <= (("@"-"@")<<11) | 0;
		m[33] <= (("@"-"@")<<11) | 64;
		m[34] <= (("@"-"@")<<11) | 48;
		m[35] <= (("@"-"@")<<11) | 10;
		m[36] <= (("@"-"@")<<11) | 1;
		m[37] <= (("@"-"@")<<11) | 0;
	end
endmodule
